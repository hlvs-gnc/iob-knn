`define KNN_ADDR_W 8  //address width
`define KNN_WDATA_W 32 //write data width
`ifndef DATA_W
 `define DATA_W 32      //cpu data width
`endif
`ifndef NBR_KNN
 `define NBR_KNN 4
`endif
`ifndef NBR_TESTP
 `define NBR_TESTP 4
`endif
